

module clk_mux (
    input       clk0_p,
    input       clk0_n,
    input       clk1_p,
    input       clk1_n,
    input       clk2,

    input [1:0] sel,

    output      clk_muxed
);

endmodule
