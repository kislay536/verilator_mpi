
 module pll_top ( 
   output clk_locked,
   output clk_out,

   input ref_clk,
   input rst,
   input bypass_en,
   input [4:0] rangeA
);


endmodule
